module IR_decoder(
input logic [31:0] ;
output logic [15:0] to_mux;
);

endmodule
