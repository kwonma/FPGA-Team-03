module top(
  input logic [1:0] key,
  input logic ir,
  input logic [7:0] but,
  output logic [2:0] snes_out);
